/* module modulo ( a, b, c);
  input [3:0] a;
  input [3:0] b;
  output reg c;
  always @(a or b) begin
    c = a % b;
  end
endmodule */